/home/patrick/wrk/proj/mcht/mcht_demo/rtl/mcht_trx.sv